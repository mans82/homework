** Profile: "SCHEMATIC1-I_sc"  [ c:\users\amir and amin\desktop\elec_finalproject\soal2_right\i_sc\i_sc-schematic1-i_sc.sim ] 

** Creating circuit file "i_sc-schematic1-i_sc.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\i_sc-SCHEMATIC1.net" 


.END
