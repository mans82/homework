** Profile: "SCHEMATIC1-Q2_LL"  [ C:\USERS\AMIR AND AMIN\DESKTOP\Elec_FinalProject\Soal2_left\soal2_left-SCHEMATIC1-Q2_LL.sim ] 

** Creating circuit file "soal2_left-SCHEMATIC1-Q2_LL.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal2_left-SCHEMATIC1.net" 


.END
