** Profile: "SCHEMATIC1-Sim"  [ e:\eec simulations\hw01s\q2\eec-hw03-q2-SCHEMATIC1-Sim.sim ] 

** Creating circuit file "eec-hw03-q2-SCHEMATIC1-Sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\eec-hw03-q2-SCHEMATIC1.net" 


.END
