** Profile: "SCHEMATIC1-mysim"  [ E:\EEC Simulations\Project\Q1\Eq2\eec - project - q1 - eq2-SCHEMATIC1-mysim.sim ] 

** Creating circuit file "eec - project - q1 - eq2-SCHEMATIC1-mysim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\eec - project - q1 - eq2-SCHEMATIC1.net" 


.END
