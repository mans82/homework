** Profile: "SCHEMATIC1-x"  [ C:\Users\Amir and Amin\Desktop\Elec_FinalProject\Soal3\soal3-SCHEMATIC1-x.sim ] 

** Creating circuit file "soal3-SCHEMATIC1-x.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 0.001 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal3-SCHEMATIC1.net" 


.END
